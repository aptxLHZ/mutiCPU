// asm file name: sra.o
module instr_rom(
    input  logic clk, rst_n,
    input  logic [13:0] i_addr,
    output logic [31:0] o_data
);
    localparam  INSTR_CNT = 12'd369;
    
    wire [0:INSTR_CNT-1] [31:0] instr_rom_cell = {
        32'h800000b7,    //0x00000000
        32'h00000113,    //0x00000004
        32'h4020df33,    //0x00000008
        32'h80000eb7,    //0x0000000c
        32'h00200193,    //0x00000010
        32'h59df1463,    //0x00000014
        32'h800000b7,    //0x00000018
        32'h00100113,    //0x0000001c
        32'h4020df33,    //0x00000020
        32'hc0000eb7,    //0x00000024
        32'h00300193,    //0x00000028
        32'h57df1863,    //0x0000002c
        32'h800000b7,    //0x00000030
        32'h00700113,    //0x00000034
        32'h4020df33,    //0x00000038
        32'hff000eb7,    //0x0000003c
        32'h00400193,    //0x00000040
        32'h55df1c63,    //0x00000044
        32'h800000b7,    //0x00000048
        32'h00e00113,    //0x0000004c
        32'h4020df33,    //0x00000050
        32'hfffe0eb7,    //0x00000054
        32'h00500193,    //0x00000058
        32'h55df1063,    //0x0000005c
        32'h800000b7,    //0x00000060
        32'h00108093,    //0x00000064
        32'h01f00113,    //0x00000068
        32'h4020df33,    //0x0000006c
        32'hfff00e93,    //0x00000070
        32'h00600193,    //0x00000074
        32'h53df1263,    //0x00000078
        32'h800000b7,    //0x0000007c
        32'hfff08093,    //0x00000080
        32'h00000113,    //0x00000084
        32'h4020df33,    //0x00000088
        32'h80000eb7,    //0x0000008c
        32'hfffe8e93,    //0x00000090
        32'h00700193,    //0x00000094
        32'h51df1263,    //0x00000098
        32'h800000b7,    //0x0000009c
        32'hfff08093,    //0x000000a0
        32'h00100113,    //0x000000a4
        32'h4020df33,    //0x000000a8
        32'h40000eb7,    //0x000000ac
        32'hfffe8e93,    //0x000000b0
        32'h00800193,    //0x000000b4
        32'h4fdf1263,    //0x000000b8
        32'h800000b7,    //0x000000bc
        32'hfff08093,    //0x000000c0
        32'h00700113,    //0x000000c4
        32'h4020df33,    //0x000000c8
        32'h01000eb7,    //0x000000cc
        32'hfffe8e93,    //0x000000d0
        32'h00900193,    //0x000000d4
        32'h4ddf1263,    //0x000000d8
        32'h800000b7,    //0x000000dc
        32'hfff08093,    //0x000000e0
        32'h00e00113,    //0x000000e4
        32'h4020df33,    //0x000000e8
        32'h00020eb7,    //0x000000ec
        32'hfffe8e93,    //0x000000f0
        32'h00a00193,    //0x000000f4
        32'h4bdf1263,    //0x000000f8
        32'h800000b7,    //0x000000fc
        32'hfff08093,    //0x00000100
        32'h01f00113,    //0x00000104
        32'h4020df33,    //0x00000108
        32'h00000e93,    //0x0000010c
        32'h00b00193,    //0x00000110
        32'h49df1463,    //0x00000114
        32'h818180b7,    //0x00000118
        32'h18108093,    //0x0000011c
        32'h00000113,    //0x00000120
        32'h4020df33,    //0x00000124
        32'h81818eb7,    //0x00000128
        32'h181e8e93,    //0x0000012c
        32'h00c00193,    //0x00000130
        32'h47df1463,    //0x00000134
        32'h818180b7,    //0x00000138
        32'h18108093,    //0x0000013c
        32'h00100113,    //0x00000140
        32'h4020df33,    //0x00000144
        32'hc0c0ceb7,    //0x00000148
        32'h0c0e8e93,    //0x0000014c
        32'h00d00193,    //0x00000150
        32'h45df1463,    //0x00000154
        32'h818180b7,    //0x00000158
        32'h18108093,    //0x0000015c
        32'h00700113,    //0x00000160
        32'h4020df33,    //0x00000164
        32'hff030eb7,    //0x00000168
        32'h303e8e93,    //0x0000016c
        32'h00e00193,    //0x00000170
        32'h43df1463,    //0x00000174
        32'h818180b7,    //0x00000178
        32'h18108093,    //0x0000017c
        32'h00e00113,    //0x00000180
        32'h4020df33,    //0x00000184
        32'hfffe0eb7,    //0x00000188
        32'h606e8e93,    //0x0000018c
        32'h00f00193,    //0x00000190
        32'h41df1463,    //0x00000194
        32'h818180b7,    //0x00000198
        32'h18108093,    //0x0000019c
        32'h01f00113,    //0x000001a0
        32'h4020df33,    //0x000001a4
        32'hfff00e93,    //0x000001a8
        32'h01000193,    //0x000001ac
        32'h3fdf1663,    //0x000001b0
        32'h818180b7,    //0x000001b4
        32'h18108093,    //0x000001b8
        32'hfc000113,    //0x000001bc
        32'h4020df33,    //0x000001c0
        32'h81818eb7,    //0x000001c4
        32'h181e8e93,    //0x000001c8
        32'h01100193,    //0x000001cc
        32'h3ddf1663,    //0x000001d0
        32'h818180b7,    //0x000001d4
        32'h18108093,    //0x000001d8
        32'hfc100113,    //0x000001dc
        32'h4020df33,    //0x000001e0
        32'hc0c0ceb7,    //0x000001e4
        32'h0c0e8e93,    //0x000001e8
        32'h01200193,    //0x000001ec
        32'h3bdf1663,    //0x000001f0
        32'h818180b7,    //0x000001f4
        32'h18108093,    //0x000001f8
        32'hfc700113,    //0x000001fc
        32'h4020df33,    //0x00000200
        32'hff030eb7,    //0x00000204
        32'h303e8e93,    //0x00000208
        32'h01300193,    //0x0000020c
        32'h39df1663,    //0x00000210
        32'h818180b7,    //0x00000214
        32'h18108093,    //0x00000218
        32'hfce00113,    //0x0000021c
        32'h4020df33,    //0x00000220
        32'hfffe0eb7,    //0x00000224
        32'h606e8e93,    //0x00000228
        32'h01400193,    //0x0000022c
        32'h37df1663,    //0x00000230
        32'h818180b7,    //0x00000234
        32'h18108093,    //0x00000238
        32'hfff00113,    //0x0000023c
        32'h4020df33,    //0x00000240
        32'hfff00e93,    //0x00000244
        32'h01500193,    //0x00000248
        32'h35df1863,    //0x0000024c
        32'h800000b7,    //0x00000250
        32'h00700113,    //0x00000254
        32'h4020d0b3,    //0x00000258
        32'hff000eb7,    //0x0000025c
        32'h01600193,    //0x00000260
        32'h33d09c63,    //0x00000264
        32'h800000b7,    //0x00000268
        32'h00e00113,    //0x0000026c
        32'h4020d133,    //0x00000270
        32'hfffe0eb7,    //0x00000274
        32'h01700193,    //0x00000278
        32'h33d11063,    //0x0000027c
        32'h00700093,    //0x00000280
        32'h4010d0b3,    //0x00000284
        32'h00000e93,    //0x00000288
        32'h01800193,    //0x0000028c
        32'h31d09663,    //0x00000290
        32'h00000213,    //0x00000294
        32'h800000b7,    //0x00000298
        32'h00700113,    //0x0000029c
        32'h4020df33,    //0x000002a0
        32'h000f0313,    //0x000002a4
        32'h00120213,    //0x000002a8
        32'h00200293,    //0x000002ac
        32'hfe5214e3,    //0x000002b0
        32'hff000eb7,    //0x000002b4
        32'h01900193,    //0x000002b8
        32'h2fd31063,    //0x000002bc
        32'h00000213,    //0x000002c0
        32'h800000b7,    //0x000002c4
        32'h00e00113,    //0x000002c8
        32'h4020df33,    //0x000002cc
        32'h00000013,    //0x000002d0
        32'h000f0313,    //0x000002d4
        32'h00120213,    //0x000002d8
        32'h00200293,    //0x000002dc
        32'hfe5212e3,    //0x000002e0
        32'hfffe0eb7,    //0x000002e4
        32'h01a00193,    //0x000002e8
        32'h2bd31863,    //0x000002ec
        32'h00000213,    //0x000002f0
        32'h800000b7,    //0x000002f4
        32'h01f00113,    //0x000002f8
        32'h4020df33,    //0x000002fc
        32'h00000013,    //0x00000300
        32'h00000013,    //0x00000304
        32'h000f0313,    //0x00000308
        32'h00120213,    //0x0000030c
        32'h00200293,    //0x00000310
        32'hfe5210e3,    //0x00000314
        32'hfff00e93,    //0x00000318
        32'h01b00193,    //0x0000031c
        32'h27d31e63,    //0x00000320
        32'h00000213,    //0x00000324
        32'h800000b7,    //0x00000328
        32'h00700113,    //0x0000032c
        32'h4020df33,    //0x00000330
        32'h00120213,    //0x00000334
        32'h00200293,    //0x00000338
        32'hfe5216e3,    //0x0000033c
        32'hff000eb7,    //0x00000340
        32'h01c00193,    //0x00000344
        32'h25df1a63,    //0x00000348
        32'h00000213,    //0x0000034c
        32'h800000b7,    //0x00000350
        32'h00e00113,    //0x00000354
        32'h00000013,    //0x00000358
        32'h4020df33,    //0x0000035c
        32'h00120213,    //0x00000360
        32'h00200293,    //0x00000364
        32'hfe5214e3,    //0x00000368
        32'hfffe0eb7,    //0x0000036c
        32'h01d00193,    //0x00000370
        32'h23df1463,    //0x00000374
        32'h00000213,    //0x00000378
        32'h800000b7,    //0x0000037c
        32'h01f00113,    //0x00000380
        32'h00000013,    //0x00000384
        32'h00000013,    //0x00000388
        32'h4020df33,    //0x0000038c
        32'h00120213,    //0x00000390
        32'h00200293,    //0x00000394
        32'hfe5212e3,    //0x00000398
        32'hfff00e93,    //0x0000039c
        32'h01e00193,    //0x000003a0
        32'h1fdf1c63,    //0x000003a4
        32'h00000213,    //0x000003a8
        32'h800000b7,    //0x000003ac
        32'h00000013,    //0x000003b0
        32'h00700113,    //0x000003b4
        32'h4020df33,    //0x000003b8
        32'h00120213,    //0x000003bc
        32'h00200293,    //0x000003c0
        32'hfe5214e3,    //0x000003c4
        32'hff000eb7,    //0x000003c8
        32'h01f00193,    //0x000003cc
        32'h1ddf1663,    //0x000003d0
        32'h00000213,    //0x000003d4
        32'h800000b7,    //0x000003d8
        32'h00000013,    //0x000003dc
        32'h00e00113,    //0x000003e0
        32'h00000013,    //0x000003e4
        32'h4020df33,    //0x000003e8
        32'h00120213,    //0x000003ec
        32'h00200293,    //0x000003f0
        32'hfe5212e3,    //0x000003f4
        32'hfffe0eb7,    //0x000003f8
        32'h02000193,    //0x000003fc
        32'h19df1e63,    //0x00000400
        32'h00000213,    //0x00000404
        32'h800000b7,    //0x00000408
        32'h00000013,    //0x0000040c
        32'h00000013,    //0x00000410
        32'h01f00113,    //0x00000414
        32'h4020df33,    //0x00000418
        32'h00120213,    //0x0000041c
        32'h00200293,    //0x00000420
        32'hfe5212e3,    //0x00000424
        32'hfff00e93,    //0x00000428
        32'h02100193,    //0x0000042c
        32'h17df1663,    //0x00000430
        32'h00000213,    //0x00000434
        32'h00700113,    //0x00000438
        32'h800000b7,    //0x0000043c
        32'h4020df33,    //0x00000440
        32'h00120213,    //0x00000444
        32'h00200293,    //0x00000448
        32'hfe5216e3,    //0x0000044c
        32'hff000eb7,    //0x00000450
        32'h02200193,    //0x00000454
        32'h15df1263,    //0x00000458
        32'h00000213,    //0x0000045c
        32'h00e00113,    //0x00000460
        32'h800000b7,    //0x00000464
        32'h00000013,    //0x00000468
        32'h4020df33,    //0x0000046c
        32'h00120213,    //0x00000470
        32'h00200293,    //0x00000474
        32'hfe5214e3,    //0x00000478
        32'hfffe0eb7,    //0x0000047c
        32'h02300193,    //0x00000480
        32'h11df1c63,    //0x00000484
        32'h00000213,    //0x00000488
        32'h01f00113,    //0x0000048c
        32'h800000b7,    //0x00000490
        32'h00000013,    //0x00000494
        32'h00000013,    //0x00000498
        32'h4020df33,    //0x0000049c
        32'h00120213,    //0x000004a0
        32'h00200293,    //0x000004a4
        32'hfe5212e3,    //0x000004a8
        32'hfff00e93,    //0x000004ac
        32'h02400193,    //0x000004b0
        32'h0fdf1463,    //0x000004b4
        32'h00000213,    //0x000004b8
        32'h00700113,    //0x000004bc
        32'h00000013,    //0x000004c0
        32'h800000b7,    //0x000004c4
        32'h4020df33,    //0x000004c8
        32'h00120213,    //0x000004cc
        32'h00200293,    //0x000004d0
        32'hfe5214e3,    //0x000004d4
        32'hff000eb7,    //0x000004d8
        32'h02500193,    //0x000004dc
        32'h0bdf1e63,    //0x000004e0
        32'h00000213,    //0x000004e4
        32'h00e00113,    //0x000004e8
        32'h00000013,    //0x000004ec
        32'h800000b7,    //0x000004f0
        32'h00000013,    //0x000004f4
        32'h4020df33,    //0x000004f8
        32'h00120213,    //0x000004fc
        32'h00200293,    //0x00000500
        32'hfe5212e3,    //0x00000504
        32'hfffe0eb7,    //0x00000508
        32'h02600193,    //0x0000050c
        32'h09df1663,    //0x00000510
        32'h00000213,    //0x00000514
        32'h01f00113,    //0x00000518
        32'h00000013,    //0x0000051c
        32'h00000013,    //0x00000520
        32'h800000b7,    //0x00000524
        32'h4020df33,    //0x00000528
        32'h00120213,    //0x0000052c
        32'h00200293,    //0x00000530
        32'hfe5212e3,    //0x00000534
        32'hfff00e93,    //0x00000538
        32'h02700193,    //0x0000053c
        32'h05df1e63,    //0x00000540
        32'h00f00093,    //0x00000544
        32'h40105133,    //0x00000548
        32'h00000e93,    //0x0000054c
        32'h02800193,    //0x00000550
        32'h05d11463,    //0x00000554
        32'h02000093,    //0x00000558
        32'h4000d133,    //0x0000055c
        32'h02000e93,    //0x00000560
        32'h02900193,    //0x00000564
        32'h03d11a63,    //0x00000568
        32'h400050b3,    //0x0000056c
        32'h00000e93,    //0x00000570
        32'h02a00193,    //0x00000574
        32'h03d09263,    //0x00000578
        32'h40000093,    //0x0000057c
        32'h00001137,    //0x00000580
        32'h80010113,    //0x00000584
        32'h4020d033,    //0x00000588
        32'h00000e93,    //0x0000058c
        32'h02b00193,    //0x00000590
        32'h01d01463,    //0x00000594
        32'h00301863,    //0x00000598
        32'h00100793,    //0x0000059c
        32'h00000213,    //0x000005a0
        32'h00320233,    //0x000005a4
        32'h00100193,    //0x000005a8
        32'h40f181b3,    //0x000005ac
        32'hc0001073,    //0x000005b0
        32'h00000000,    //0x000005b4
        32'h00000000,    //0x000005b8
        32'h00000000,    //0x000005bc
        32'h00000000    //0x000005c0
    };
    
    logic [11:0] instr_index;
    logic [31:0] data;
    
    assign instr_index = i_addr[13:2];
    assign data = (instr_index>=INSTR_CNT) ? 0 : instr_rom_cell[instr_index];
    
    always @ (posedge clk or negedge rst_n)
        if(~rst_n)
            o_data <= 0;
        else
            o_data <= data;

endmodule
