// asm file name: lbu.o
module instr_rom(
    input  logic clk, rst_n,
    input  logic [13:0] i_addr,
    output logic [31:0] o_data
);
    localparam  INSTR_CNT = 12'd1205;
    
    wire [0:INSTR_CNT-1] [31:0] instr_rom_cell = {
        32'h00001097,    //0x00000000
        32'h26c08093,    //0x00000004
        32'h0000cf03,    //0x00000008
        32'h0ff00e93,    //0x0000000c
        32'h00200193,    //0x00000010
        32'h23df1c63,    //0x00000014
        32'h00001097,    //0x00000018
        32'h25408093,    //0x0000001c
        32'h0010cf03,    //0x00000020
        32'h00000e93,    //0x00000024
        32'h00300193,    //0x00000028
        32'h23df1063,    //0x0000002c
        32'h00001097,    //0x00000030
        32'h23c08093,    //0x00000034
        32'h0020cf03,    //0x00000038
        32'h0f000e93,    //0x0000003c
        32'h00400193,    //0x00000040
        32'h21df1463,    //0x00000044
        32'h00001097,    //0x00000048
        32'h22408093,    //0x0000004c
        32'h0030cf03,    //0x00000050
        32'h00f00e93,    //0x00000054
        32'h00500193,    //0x00000058
        32'h1fdf1863,    //0x0000005c
        32'h00001097,    //0x00000060
        32'h20f08093,    //0x00000064
        32'hffd0cf03,    //0x00000068
        32'h0ff00e93,    //0x0000006c
        32'h00600193,    //0x00000070
        32'h1ddf1c63,    //0x00000074
        32'h00001097,    //0x00000078
        32'h1f708093,    //0x0000007c
        32'hffe0cf03,    //0x00000080
        32'h00000e93,    //0x00000084
        32'h00700193,    //0x00000088
        32'h1ddf1063,    //0x0000008c
        32'h00001097,    //0x00000090
        32'h1df08093,    //0x00000094
        32'hfff0cf03,    //0x00000098
        32'h0f000e93,    //0x0000009c
        32'h00800193,    //0x000000a0
        32'h1bdf1463,    //0x000000a4
        32'h00001097,    //0x000000a8
        32'h1c708093,    //0x000000ac
        32'h0000cf03,    //0x000000b0
        32'h00f00e93,    //0x000000b4
        32'h00900193,    //0x000000b8
        32'h19df1863,    //0x000000bc
        32'h00001097,    //0x000000c0
        32'h1ac08093,    //0x000000c4
        32'hfe008093,    //0x000000c8
        32'h0200c283,    //0x000000cc
        32'h0ff00e93,    //0x000000d0
        32'h00a00193,    //0x000000d4
        32'h17d29a63,    //0x000000d8
        32'h00001097,    //0x000000dc
        32'h19008093,    //0x000000e0
        32'hffa08093,    //0x000000e4
        32'h0070c283,    //0x000000e8
        32'h00000e93,    //0x000000ec
        32'h00b00193,    //0x000000f0
        32'h15d29c63,    //0x000000f4
        32'h00c00193,    //0x000000f8
        32'h00000213,    //0x000000fc
        32'h00001097,    //0x00000100
        32'h16d08093,    //0x00000104
        32'h0010cf03,    //0x00000108
        32'h000f0313,    //0x0000010c
        32'h0f000e93,    //0x00000110
        32'h13d31c63,    //0x00000114
        32'h00120213,    //0x00000118
        32'h00200293,    //0x0000011c
        32'hfe5210e3,    //0x00000120
        32'h00d00193,    //0x00000124
        32'h00000213,    //0x00000128
        32'h00001097,    //0x0000012c
        32'h14208093,    //0x00000130
        32'h0010cf03,    //0x00000134
        32'h00000013,    //0x00000138
        32'h000f0313,    //0x0000013c
        32'h00f00e93,    //0x00000140
        32'h11d31463,    //0x00000144
        32'h00120213,    //0x00000148
        32'h00200293,    //0x0000014c
        32'hfc521ee3,    //0x00000150
        32'h00e00193,    //0x00000154
        32'h00000213,    //0x00000158
        32'h00001097,    //0x0000015c
        32'h11008093,    //0x00000160
        32'h0010cf03,    //0x00000164
        32'h00000013,    //0x00000168
        32'h00000013,    //0x0000016c
        32'h000f0313,    //0x00000170
        32'h00000e93,    //0x00000174
        32'h0dd31a63,    //0x00000178
        32'h00120213,    //0x0000017c
        32'h00200293,    //0x00000180
        32'hfc521ce3,    //0x00000184
        32'h00f00193,    //0x00000188
        32'h00000213,    //0x0000018c
        32'h00001097,    //0x00000190
        32'h0dd08093,    //0x00000194
        32'h0010cf03,    //0x00000198
        32'h0f000e93,    //0x0000019c
        32'h0bdf1663,    //0x000001a0
        32'h00120213,    //0x000001a4
        32'h00200293,    //0x000001a8
        32'hfe5212e3,    //0x000001ac
        32'h01000193,    //0x000001b0
        32'h00000213,    //0x000001b4
        32'h00001097,    //0x000001b8
        32'h0b608093,    //0x000001bc
        32'h00000013,    //0x000001c0
        32'h0010cf03,    //0x000001c4
        32'h00f00e93,    //0x000001c8
        32'h09df1063,    //0x000001cc
        32'h00120213,    //0x000001d0
        32'h00200293,    //0x000001d4
        32'hfe5210e3,    //0x000001d8
        32'h01100193,    //0x000001dc
        32'h00000213,    //0x000001e0
        32'h00001097,    //0x000001e4
        32'h08808093,    //0x000001e8
        32'h00000013,    //0x000001ec
        32'h00000013,    //0x000001f0
        32'h0010cf03,    //0x000001f4
        32'h00000e93,    //0x000001f8
        32'h05df1863,    //0x000001fc
        32'h00120213,    //0x00000200
        32'h00200293,    //0x00000204
        32'hfc521ee3,    //0x00000208
        32'h00001297,    //0x0000020c
        32'h06028293,    //0x00000210
        32'h0002c103,    //0x00000214
        32'h00200113,    //0x00000218
        32'h00200e93,    //0x0000021c
        32'h01200193,    //0x00000220
        32'h03d11463,    //0x00000224
        32'h00001297,    //0x00000228
        32'h04428293,    //0x0000022c
        32'h0002c103,    //0x00000230
        32'h00000013,    //0x00000234
        32'h00200113,    //0x00000238
        32'h00200e93,    //0x0000023c
        32'h01300193,    //0x00000240
        32'h01d11463,    //0x00000244
        32'h00301863,    //0x00000248
        32'h00100793,    //0x0000024c
        32'h00000213,    //0x00000250
        32'h00320233,    //0x00000254
        32'h00100193,    //0x00000258
        32'h40f181b3,    //0x0000025c
        32'hc0001073,    //0x00000260
        32'h00000000,    //0x00000264
        32'h00000000,    //0x00000268
        32'h00000000,    //0x0000026c
        32'h00000000,    //0x00000270
        32'h00000000,    //0x00000274
        32'h00000000,    //0x00000278
        32'h00000000,    //0x0000027c
        32'h00000000,    //0x00000280
        32'h00000000,    //0x00000284
        32'h00000000,    //0x00000288
        32'h00000000,    //0x0000028c
        32'h00000000,    //0x00000290
        32'h00000000,    //0x00000294
        32'h00000000,    //0x00000298
        32'h00000000,    //0x0000029c
        32'h00000000,    //0x000002a0
        32'h00000000,    //0x000002a4
        32'h00000000,    //0x000002a8
        32'h00000000,    //0x000002ac
        32'h00000000,    //0x000002b0
        32'h00000000,    //0x000002b4
        32'h00000000,    //0x000002b8
        32'h00000000,    //0x000002bc
        32'h00000000,    //0x000002c0
        32'h00000000,    //0x000002c4
        32'h00000000,    //0x000002c8
        32'h00000000,    //0x000002cc
        32'h00000000,    //0x000002d0
        32'h00000000,    //0x000002d4
        32'h00000000,    //0x000002d8
        32'h00000000,    //0x000002dc
        32'h00000000,    //0x000002e0
        32'h00000000,    //0x000002e4
        32'h00000000,    //0x000002e8
        32'h00000000,    //0x000002ec
        32'h00000000,    //0x000002f0
        32'h00000000,    //0x000002f4
        32'h00000000,    //0x000002f8
        32'h00000000,    //0x000002fc
        32'h00000000,    //0x00000300
        32'h00000000,    //0x00000304
        32'h00000000,    //0x00000308
        32'h00000000,    //0x0000030c
        32'h00000000,    //0x00000310
        32'h00000000,    //0x00000314
        32'h00000000,    //0x00000318
        32'h00000000,    //0x0000031c
        32'h00000000,    //0x00000320
        32'h00000000,    //0x00000324
        32'h00000000,    //0x00000328
        32'h00000000,    //0x0000032c
        32'h00000000,    //0x00000330
        32'h00000000,    //0x00000334
        32'h00000000,    //0x00000338
        32'h00000000,    //0x0000033c
        32'h00000000,    //0x00000340
        32'h00000000,    //0x00000344
        32'h00000000,    //0x00000348
        32'h00000000,    //0x0000034c
        32'h00000000,    //0x00000350
        32'h00000000,    //0x00000354
        32'h00000000,    //0x00000358
        32'h00000000,    //0x0000035c
        32'h00000000,    //0x00000360
        32'h00000000,    //0x00000364
        32'h00000000,    //0x00000368
        32'h00000000,    //0x0000036c
        32'h00000000,    //0x00000370
        32'h00000000,    //0x00000374
        32'h00000000,    //0x00000378
        32'h00000000,    //0x0000037c
        32'h00000000,    //0x00000380
        32'h00000000,    //0x00000384
        32'h00000000,    //0x00000388
        32'h00000000,    //0x0000038c
        32'h00000000,    //0x00000390
        32'h00000000,    //0x00000394
        32'h00000000,    //0x00000398
        32'h00000000,    //0x0000039c
        32'h00000000,    //0x000003a0
        32'h00000000,    //0x000003a4
        32'h00000000,    //0x000003a8
        32'h00000000,    //0x000003ac
        32'h00000000,    //0x000003b0
        32'h00000000,    //0x000003b4
        32'h00000000,    //0x000003b8
        32'h00000000,    //0x000003bc
        32'h00000000,    //0x000003c0
        32'h00000000,    //0x000003c4
        32'h00000000,    //0x000003c8
        32'h00000000,    //0x000003cc
        32'h00000000,    //0x000003d0
        32'h00000000,    //0x000003d4
        32'h00000000,    //0x000003d8
        32'h00000000,    //0x000003dc
        32'h00000000,    //0x000003e0
        32'h00000000,    //0x000003e4
        32'h00000000,    //0x000003e8
        32'h00000000,    //0x000003ec
        32'h00000000,    //0x000003f0
        32'h00000000,    //0x000003f4
        32'h00000000,    //0x000003f8
        32'h00000000,    //0x000003fc
        32'h00000000,    //0x00000400
        32'h00000000,    //0x00000404
        32'h00000000,    //0x00000408
        32'h00000000,    //0x0000040c
        32'h00000000,    //0x00000410
        32'h00000000,    //0x00000414
        32'h00000000,    //0x00000418
        32'h00000000,    //0x0000041c
        32'h00000000,    //0x00000420
        32'h00000000,    //0x00000424
        32'h00000000,    //0x00000428
        32'h00000000,    //0x0000042c
        32'h00000000,    //0x00000430
        32'h00000000,    //0x00000434
        32'h00000000,    //0x00000438
        32'h00000000,    //0x0000043c
        32'h00000000,    //0x00000440
        32'h00000000,    //0x00000444
        32'h00000000,    //0x00000448
        32'h00000000,    //0x0000044c
        32'h00000000,    //0x00000450
        32'h00000000,    //0x00000454
        32'h00000000,    //0x00000458
        32'h00000000,    //0x0000045c
        32'h00000000,    //0x00000460
        32'h00000000,    //0x00000464
        32'h00000000,    //0x00000468
        32'h00000000,    //0x0000046c
        32'h00000000,    //0x00000470
        32'h00000000,    //0x00000474
        32'h00000000,    //0x00000478
        32'h00000000,    //0x0000047c
        32'h00000000,    //0x00000480
        32'h00000000,    //0x00000484
        32'h00000000,    //0x00000488
        32'h00000000,    //0x0000048c
        32'h00000000,    //0x00000490
        32'h00000000,    //0x00000494
        32'h00000000,    //0x00000498
        32'h00000000,    //0x0000049c
        32'h00000000,    //0x000004a0
        32'h00000000,    //0x000004a4
        32'h00000000,    //0x000004a8
        32'h00000000,    //0x000004ac
        32'h00000000,    //0x000004b0
        32'h00000000,    //0x000004b4
        32'h00000000,    //0x000004b8
        32'h00000000,    //0x000004bc
        32'h00000000,    //0x000004c0
        32'h00000000,    //0x000004c4
        32'h00000000,    //0x000004c8
        32'h00000000,    //0x000004cc
        32'h00000000,    //0x000004d0
        32'h00000000,    //0x000004d4
        32'h00000000,    //0x000004d8
        32'h00000000,    //0x000004dc
        32'h00000000,    //0x000004e0
        32'h00000000,    //0x000004e4
        32'h00000000,    //0x000004e8
        32'h00000000,    //0x000004ec
        32'h00000000,    //0x000004f0
        32'h00000000,    //0x000004f4
        32'h00000000,    //0x000004f8
        32'h00000000,    //0x000004fc
        32'h00000000,    //0x00000500
        32'h00000000,    //0x00000504
        32'h00000000,    //0x00000508
        32'h00000000,    //0x0000050c
        32'h00000000,    //0x00000510
        32'h00000000,    //0x00000514
        32'h00000000,    //0x00000518
        32'h00000000,    //0x0000051c
        32'h00000000,    //0x00000520
        32'h00000000,    //0x00000524
        32'h00000000,    //0x00000528
        32'h00000000,    //0x0000052c
        32'h00000000,    //0x00000530
        32'h00000000,    //0x00000534
        32'h00000000,    //0x00000538
        32'h00000000,    //0x0000053c
        32'h00000000,    //0x00000540
        32'h00000000,    //0x00000544
        32'h00000000,    //0x00000548
        32'h00000000,    //0x0000054c
        32'h00000000,    //0x00000550
        32'h00000000,    //0x00000554
        32'h00000000,    //0x00000558
        32'h00000000,    //0x0000055c
        32'h00000000,    //0x00000560
        32'h00000000,    //0x00000564
        32'h00000000,    //0x00000568
        32'h00000000,    //0x0000056c
        32'h00000000,    //0x00000570
        32'h00000000,    //0x00000574
        32'h00000000,    //0x00000578
        32'h00000000,    //0x0000057c
        32'h00000000,    //0x00000580
        32'h00000000,    //0x00000584
        32'h00000000,    //0x00000588
        32'h00000000,    //0x0000058c
        32'h00000000,    //0x00000590
        32'h00000000,    //0x00000594
        32'h00000000,    //0x00000598
        32'h00000000,    //0x0000059c
        32'h00000000,    //0x000005a0
        32'h00000000,    //0x000005a4
        32'h00000000,    //0x000005a8
        32'h00000000,    //0x000005ac
        32'h00000000,    //0x000005b0
        32'h00000000,    //0x000005b4
        32'h00000000,    //0x000005b8
        32'h00000000,    //0x000005bc
        32'h00000000,    //0x000005c0
        32'h00000000,    //0x000005c4
        32'h00000000,    //0x000005c8
        32'h00000000,    //0x000005cc
        32'h00000000,    //0x000005d0
        32'h00000000,    //0x000005d4
        32'h00000000,    //0x000005d8
        32'h00000000,    //0x000005dc
        32'h00000000,    //0x000005e0
        32'h00000000,    //0x000005e4
        32'h00000000,    //0x000005e8
        32'h00000000,    //0x000005ec
        32'h00000000,    //0x000005f0
        32'h00000000,    //0x000005f4
        32'h00000000,    //0x000005f8
        32'h00000000,    //0x000005fc
        32'h00000000,    //0x00000600
        32'h00000000,    //0x00000604
        32'h00000000,    //0x00000608
        32'h00000000,    //0x0000060c
        32'h00000000,    //0x00000610
        32'h00000000,    //0x00000614
        32'h00000000,    //0x00000618
        32'h00000000,    //0x0000061c
        32'h00000000,    //0x00000620
        32'h00000000,    //0x00000624
        32'h00000000,    //0x00000628
        32'h00000000,    //0x0000062c
        32'h00000000,    //0x00000630
        32'h00000000,    //0x00000634
        32'h00000000,    //0x00000638
        32'h00000000,    //0x0000063c
        32'h00000000,    //0x00000640
        32'h00000000,    //0x00000644
        32'h00000000,    //0x00000648
        32'h00000000,    //0x0000064c
        32'h00000000,    //0x00000650
        32'h00000000,    //0x00000654
        32'h00000000,    //0x00000658
        32'h00000000,    //0x0000065c
        32'h00000000,    //0x00000660
        32'h00000000,    //0x00000664
        32'h00000000,    //0x00000668
        32'h00000000,    //0x0000066c
        32'h00000000,    //0x00000670
        32'h00000000,    //0x00000674
        32'h00000000,    //0x00000678
        32'h00000000,    //0x0000067c
        32'h00000000,    //0x00000680
        32'h00000000,    //0x00000684
        32'h00000000,    //0x00000688
        32'h00000000,    //0x0000068c
        32'h00000000,    //0x00000690
        32'h00000000,    //0x00000694
        32'h00000000,    //0x00000698
        32'h00000000,    //0x0000069c
        32'h00000000,    //0x000006a0
        32'h00000000,    //0x000006a4
        32'h00000000,    //0x000006a8
        32'h00000000,    //0x000006ac
        32'h00000000,    //0x000006b0
        32'h00000000,    //0x000006b4
        32'h00000000,    //0x000006b8
        32'h00000000,    //0x000006bc
        32'h00000000,    //0x000006c0
        32'h00000000,    //0x000006c4
        32'h00000000,    //0x000006c8
        32'h00000000,    //0x000006cc
        32'h00000000,    //0x000006d0
        32'h00000000,    //0x000006d4
        32'h00000000,    //0x000006d8
        32'h00000000,    //0x000006dc
        32'h00000000,    //0x000006e0
        32'h00000000,    //0x000006e4
        32'h00000000,    //0x000006e8
        32'h00000000,    //0x000006ec
        32'h00000000,    //0x000006f0
        32'h00000000,    //0x000006f4
        32'h00000000,    //0x000006f8
        32'h00000000,    //0x000006fc
        32'h00000000,    //0x00000700
        32'h00000000,    //0x00000704
        32'h00000000,    //0x00000708
        32'h00000000,    //0x0000070c
        32'h00000000,    //0x00000710
        32'h00000000,    //0x00000714
        32'h00000000,    //0x00000718
        32'h00000000,    //0x0000071c
        32'h00000000,    //0x00000720
        32'h00000000,    //0x00000724
        32'h00000000,    //0x00000728
        32'h00000000,    //0x0000072c
        32'h00000000,    //0x00000730
        32'h00000000,    //0x00000734
        32'h00000000,    //0x00000738
        32'h00000000,    //0x0000073c
        32'h00000000,    //0x00000740
        32'h00000000,    //0x00000744
        32'h00000000,    //0x00000748
        32'h00000000,    //0x0000074c
        32'h00000000,    //0x00000750
        32'h00000000,    //0x00000754
        32'h00000000,    //0x00000758
        32'h00000000,    //0x0000075c
        32'h00000000,    //0x00000760
        32'h00000000,    //0x00000764
        32'h00000000,    //0x00000768
        32'h00000000,    //0x0000076c
        32'h00000000,    //0x00000770
        32'h00000000,    //0x00000774
        32'h00000000,    //0x00000778
        32'h00000000,    //0x0000077c
        32'h00000000,    //0x00000780
        32'h00000000,    //0x00000784
        32'h00000000,    //0x00000788
        32'h00000000,    //0x0000078c
        32'h00000000,    //0x00000790
        32'h00000000,    //0x00000794
        32'h00000000,    //0x00000798
        32'h00000000,    //0x0000079c
        32'h00000000,    //0x000007a0
        32'h00000000,    //0x000007a4
        32'h00000000,    //0x000007a8
        32'h00000000,    //0x000007ac
        32'h00000000,    //0x000007b0
        32'h00000000,    //0x000007b4
        32'h00000000,    //0x000007b8
        32'h00000000,    //0x000007bc
        32'h00000000,    //0x000007c0
        32'h00000000,    //0x000007c4
        32'h00000000,    //0x000007c8
        32'h00000000,    //0x000007cc
        32'h00000000,    //0x000007d0
        32'h00000000,    //0x000007d4
        32'h00000000,    //0x000007d8
        32'h00000000,    //0x000007dc
        32'h00000000,    //0x000007e0
        32'h00000000,    //0x000007e4
        32'h00000000,    //0x000007e8
        32'h00000000,    //0x000007ec
        32'h00000000,    //0x000007f0
        32'h00000000,    //0x000007f4
        32'h00000000,    //0x000007f8
        32'h00000000,    //0x000007fc
        32'h00000000,    //0x00000800
        32'h00000000,    //0x00000804
        32'h00000000,    //0x00000808
        32'h00000000,    //0x0000080c
        32'h00000000,    //0x00000810
        32'h00000000,    //0x00000814
        32'h00000000,    //0x00000818
        32'h00000000,    //0x0000081c
        32'h00000000,    //0x00000820
        32'h00000000,    //0x00000824
        32'h00000000,    //0x00000828
        32'h00000000,    //0x0000082c
        32'h00000000,    //0x00000830
        32'h00000000,    //0x00000834
        32'h00000000,    //0x00000838
        32'h00000000,    //0x0000083c
        32'h00000000,    //0x00000840
        32'h00000000,    //0x00000844
        32'h00000000,    //0x00000848
        32'h00000000,    //0x0000084c
        32'h00000000,    //0x00000850
        32'h00000000,    //0x00000854
        32'h00000000,    //0x00000858
        32'h00000000,    //0x0000085c
        32'h00000000,    //0x00000860
        32'h00000000,    //0x00000864
        32'h00000000,    //0x00000868
        32'h00000000,    //0x0000086c
        32'h00000000,    //0x00000870
        32'h00000000,    //0x00000874
        32'h00000000,    //0x00000878
        32'h00000000,    //0x0000087c
        32'h00000000,    //0x00000880
        32'h00000000,    //0x00000884
        32'h00000000,    //0x00000888
        32'h00000000,    //0x0000088c
        32'h00000000,    //0x00000890
        32'h00000000,    //0x00000894
        32'h00000000,    //0x00000898
        32'h00000000,    //0x0000089c
        32'h00000000,    //0x000008a0
        32'h00000000,    //0x000008a4
        32'h00000000,    //0x000008a8
        32'h00000000,    //0x000008ac
        32'h00000000,    //0x000008b0
        32'h00000000,    //0x000008b4
        32'h00000000,    //0x000008b8
        32'h00000000,    //0x000008bc
        32'h00000000,    //0x000008c0
        32'h00000000,    //0x000008c4
        32'h00000000,    //0x000008c8
        32'h00000000,    //0x000008cc
        32'h00000000,    //0x000008d0
        32'h00000000,    //0x000008d4
        32'h00000000,    //0x000008d8
        32'h00000000,    //0x000008dc
        32'h00000000,    //0x000008e0
        32'h00000000,    //0x000008e4
        32'h00000000,    //0x000008e8
        32'h00000000,    //0x000008ec
        32'h00000000,    //0x000008f0
        32'h00000000,    //0x000008f4
        32'h00000000,    //0x000008f8
        32'h00000000,    //0x000008fc
        32'h00000000,    //0x00000900
        32'h00000000,    //0x00000904
        32'h00000000,    //0x00000908
        32'h00000000,    //0x0000090c
        32'h00000000,    //0x00000910
        32'h00000000,    //0x00000914
        32'h00000000,    //0x00000918
        32'h00000000,    //0x0000091c
        32'h00000000,    //0x00000920
        32'h00000000,    //0x00000924
        32'h00000000,    //0x00000928
        32'h00000000,    //0x0000092c
        32'h00000000,    //0x00000930
        32'h00000000,    //0x00000934
        32'h00000000,    //0x00000938
        32'h00000000,    //0x0000093c
        32'h00000000,    //0x00000940
        32'h00000000,    //0x00000944
        32'h00000000,    //0x00000948
        32'h00000000,    //0x0000094c
        32'h00000000,    //0x00000950
        32'h00000000,    //0x00000954
        32'h00000000,    //0x00000958
        32'h00000000,    //0x0000095c
        32'h00000000,    //0x00000960
        32'h00000000,    //0x00000964
        32'h00000000,    //0x00000968
        32'h00000000,    //0x0000096c
        32'h00000000,    //0x00000970
        32'h00000000,    //0x00000974
        32'h00000000,    //0x00000978
        32'h00000000,    //0x0000097c
        32'h00000000,    //0x00000980
        32'h00000000,    //0x00000984
        32'h00000000,    //0x00000988
        32'h00000000,    //0x0000098c
        32'h00000000,    //0x00000990
        32'h00000000,    //0x00000994
        32'h00000000,    //0x00000998
        32'h00000000,    //0x0000099c
        32'h00000000,    //0x000009a0
        32'h00000000,    //0x000009a4
        32'h00000000,    //0x000009a8
        32'h00000000,    //0x000009ac
        32'h00000000,    //0x000009b0
        32'h00000000,    //0x000009b4
        32'h00000000,    //0x000009b8
        32'h00000000,    //0x000009bc
        32'h00000000,    //0x000009c0
        32'h00000000,    //0x000009c4
        32'h00000000,    //0x000009c8
        32'h00000000,    //0x000009cc
        32'h00000000,    //0x000009d0
        32'h00000000,    //0x000009d4
        32'h00000000,    //0x000009d8
        32'h00000000,    //0x000009dc
        32'h00000000,    //0x000009e0
        32'h00000000,    //0x000009e4
        32'h00000000,    //0x000009e8
        32'h00000000,    //0x000009ec
        32'h00000000,    //0x000009f0
        32'h00000000,    //0x000009f4
        32'h00000000,    //0x000009f8
        32'h00000000,    //0x000009fc
        32'h00000000,    //0x00000a00
        32'h00000000,    //0x00000a04
        32'h00000000,    //0x00000a08
        32'h00000000,    //0x00000a0c
        32'h00000000,    //0x00000a10
        32'h00000000,    //0x00000a14
        32'h00000000,    //0x00000a18
        32'h00000000,    //0x00000a1c
        32'h00000000,    //0x00000a20
        32'h00000000,    //0x00000a24
        32'h00000000,    //0x00000a28
        32'h00000000,    //0x00000a2c
        32'h00000000,    //0x00000a30
        32'h00000000,    //0x00000a34
        32'h00000000,    //0x00000a38
        32'h00000000,    //0x00000a3c
        32'h00000000,    //0x00000a40
        32'h00000000,    //0x00000a44
        32'h00000000,    //0x00000a48
        32'h00000000,    //0x00000a4c
        32'h00000000,    //0x00000a50
        32'h00000000,    //0x00000a54
        32'h00000000,    //0x00000a58
        32'h00000000,    //0x00000a5c
        32'h00000000,    //0x00000a60
        32'h00000000,    //0x00000a64
        32'h00000000,    //0x00000a68
        32'h00000000,    //0x00000a6c
        32'h00000000,    //0x00000a70
        32'h00000000,    //0x00000a74
        32'h00000000,    //0x00000a78
        32'h00000000,    //0x00000a7c
        32'h00000000,    //0x00000a80
        32'h00000000,    //0x00000a84
        32'h00000000,    //0x00000a88
        32'h00000000,    //0x00000a8c
        32'h00000000,    //0x00000a90
        32'h00000000,    //0x00000a94
        32'h00000000,    //0x00000a98
        32'h00000000,    //0x00000a9c
        32'h00000000,    //0x00000aa0
        32'h00000000,    //0x00000aa4
        32'h00000000,    //0x00000aa8
        32'h00000000,    //0x00000aac
        32'h00000000,    //0x00000ab0
        32'h00000000,    //0x00000ab4
        32'h00000000,    //0x00000ab8
        32'h00000000,    //0x00000abc
        32'h00000000,    //0x00000ac0
        32'h00000000,    //0x00000ac4
        32'h00000000,    //0x00000ac8
        32'h00000000,    //0x00000acc
        32'h00000000,    //0x00000ad0
        32'h00000000,    //0x00000ad4
        32'h00000000,    //0x00000ad8
        32'h00000000,    //0x00000adc
        32'h00000000,    //0x00000ae0
        32'h00000000,    //0x00000ae4
        32'h00000000,    //0x00000ae8
        32'h00000000,    //0x00000aec
        32'h00000000,    //0x00000af0
        32'h00000000,    //0x00000af4
        32'h00000000,    //0x00000af8
        32'h00000000,    //0x00000afc
        32'h00000000,    //0x00000b00
        32'h00000000,    //0x00000b04
        32'h00000000,    //0x00000b08
        32'h00000000,    //0x00000b0c
        32'h00000000,    //0x00000b10
        32'h00000000,    //0x00000b14
        32'h00000000,    //0x00000b18
        32'h00000000,    //0x00000b1c
        32'h00000000,    //0x00000b20
        32'h00000000,    //0x00000b24
        32'h00000000,    //0x00000b28
        32'h00000000,    //0x00000b2c
        32'h00000000,    //0x00000b30
        32'h00000000,    //0x00000b34
        32'h00000000,    //0x00000b38
        32'h00000000,    //0x00000b3c
        32'h00000000,    //0x00000b40
        32'h00000000,    //0x00000b44
        32'h00000000,    //0x00000b48
        32'h00000000,    //0x00000b4c
        32'h00000000,    //0x00000b50
        32'h00000000,    //0x00000b54
        32'h00000000,    //0x00000b58
        32'h00000000,    //0x00000b5c
        32'h00000000,    //0x00000b60
        32'h00000000,    //0x00000b64
        32'h00000000,    //0x00000b68
        32'h00000000,    //0x00000b6c
        32'h00000000,    //0x00000b70
        32'h00000000,    //0x00000b74
        32'h00000000,    //0x00000b78
        32'h00000000,    //0x00000b7c
        32'h00000000,    //0x00000b80
        32'h00000000,    //0x00000b84
        32'h00000000,    //0x00000b88
        32'h00000000,    //0x00000b8c
        32'h00000000,    //0x00000b90
        32'h00000000,    //0x00000b94
        32'h00000000,    //0x00000b98
        32'h00000000,    //0x00000b9c
        32'h00000000,    //0x00000ba0
        32'h00000000,    //0x00000ba4
        32'h00000000,    //0x00000ba8
        32'h00000000,    //0x00000bac
        32'h00000000,    //0x00000bb0
        32'h00000000,    //0x00000bb4
        32'h00000000,    //0x00000bb8
        32'h00000000,    //0x00000bbc
        32'h00000000,    //0x00000bc0
        32'h00000000,    //0x00000bc4
        32'h00000000,    //0x00000bc8
        32'h00000000,    //0x00000bcc
        32'h00000000,    //0x00000bd0
        32'h00000000,    //0x00000bd4
        32'h00000000,    //0x00000bd8
        32'h00000000,    //0x00000bdc
        32'h00000000,    //0x00000be0
        32'h00000000,    //0x00000be4
        32'h00000000,    //0x00000be8
        32'h00000000,    //0x00000bec
        32'h00000000,    //0x00000bf0
        32'h00000000,    //0x00000bf4
        32'h00000000,    //0x00000bf8
        32'h00000000,    //0x00000bfc
        32'h00000000,    //0x00000c00
        32'h00000000,    //0x00000c04
        32'h00000000,    //0x00000c08
        32'h00000000,    //0x00000c0c
        32'h00000000,    //0x00000c10
        32'h00000000,    //0x00000c14
        32'h00000000,    //0x00000c18
        32'h00000000,    //0x00000c1c
        32'h00000000,    //0x00000c20
        32'h00000000,    //0x00000c24
        32'h00000000,    //0x00000c28
        32'h00000000,    //0x00000c2c
        32'h00000000,    //0x00000c30
        32'h00000000,    //0x00000c34
        32'h00000000,    //0x00000c38
        32'h00000000,    //0x00000c3c
        32'h00000000,    //0x00000c40
        32'h00000000,    //0x00000c44
        32'h00000000,    //0x00000c48
        32'h00000000,    //0x00000c4c
        32'h00000000,    //0x00000c50
        32'h00000000,    //0x00000c54
        32'h00000000,    //0x00000c58
        32'h00000000,    //0x00000c5c
        32'h00000000,    //0x00000c60
        32'h00000000,    //0x00000c64
        32'h00000000,    //0x00000c68
        32'h00000000,    //0x00000c6c
        32'h00000000,    //0x00000c70
        32'h00000000,    //0x00000c74
        32'h00000000,    //0x00000c78
        32'h00000000,    //0x00000c7c
        32'h00000000,    //0x00000c80
        32'h00000000,    //0x00000c84
        32'h00000000,    //0x00000c88
        32'h00000000,    //0x00000c8c
        32'h00000000,    //0x00000c90
        32'h00000000,    //0x00000c94
        32'h00000000,    //0x00000c98
        32'h00000000,    //0x00000c9c
        32'h00000000,    //0x00000ca0
        32'h00000000,    //0x00000ca4
        32'h00000000,    //0x00000ca8
        32'h00000000,    //0x00000cac
        32'h00000000,    //0x00000cb0
        32'h00000000,    //0x00000cb4
        32'h00000000,    //0x00000cb8
        32'h00000000,    //0x00000cbc
        32'h00000000,    //0x00000cc0
        32'h00000000,    //0x00000cc4
        32'h00000000,    //0x00000cc8
        32'h00000000,    //0x00000ccc
        32'h00000000,    //0x00000cd0
        32'h00000000,    //0x00000cd4
        32'h00000000,    //0x00000cd8
        32'h00000000,    //0x00000cdc
        32'h00000000,    //0x00000ce0
        32'h00000000,    //0x00000ce4
        32'h00000000,    //0x00000ce8
        32'h00000000,    //0x00000cec
        32'h00000000,    //0x00000cf0
        32'h00000000,    //0x00000cf4
        32'h00000000,    //0x00000cf8
        32'h00000000,    //0x00000cfc
        32'h00000000,    //0x00000d00
        32'h00000000,    //0x00000d04
        32'h00000000,    //0x00000d08
        32'h00000000,    //0x00000d0c
        32'h00000000,    //0x00000d10
        32'h00000000,    //0x00000d14
        32'h00000000,    //0x00000d18
        32'h00000000,    //0x00000d1c
        32'h00000000,    //0x00000d20
        32'h00000000,    //0x00000d24
        32'h00000000,    //0x00000d28
        32'h00000000,    //0x00000d2c
        32'h00000000,    //0x00000d30
        32'h00000000,    //0x00000d34
        32'h00000000,    //0x00000d38
        32'h00000000,    //0x00000d3c
        32'h00000000,    //0x00000d40
        32'h00000000,    //0x00000d44
        32'h00000000,    //0x00000d48
        32'h00000000,    //0x00000d4c
        32'h00000000,    //0x00000d50
        32'h00000000,    //0x00000d54
        32'h00000000,    //0x00000d58
        32'h00000000,    //0x00000d5c
        32'h00000000,    //0x00000d60
        32'h00000000,    //0x00000d64
        32'h00000000,    //0x00000d68
        32'h00000000,    //0x00000d6c
        32'h00000000,    //0x00000d70
        32'h00000000,    //0x00000d74
        32'h00000000,    //0x00000d78
        32'h00000000,    //0x00000d7c
        32'h00000000,    //0x00000d80
        32'h00000000,    //0x00000d84
        32'h00000000,    //0x00000d88
        32'h00000000,    //0x00000d8c
        32'h00000000,    //0x00000d90
        32'h00000000,    //0x00000d94
        32'h00000000,    //0x00000d98
        32'h00000000,    //0x00000d9c
        32'h00000000,    //0x00000da0
        32'h00000000,    //0x00000da4
        32'h00000000,    //0x00000da8
        32'h00000000,    //0x00000dac
        32'h00000000,    //0x00000db0
        32'h00000000,    //0x00000db4
        32'h00000000,    //0x00000db8
        32'h00000000,    //0x00000dbc
        32'h00000000,    //0x00000dc0
        32'h00000000,    //0x00000dc4
        32'h00000000,    //0x00000dc8
        32'h00000000,    //0x00000dcc
        32'h00000000,    //0x00000dd0
        32'h00000000,    //0x00000dd4
        32'h00000000,    //0x00000dd8
        32'h00000000,    //0x00000ddc
        32'h00000000,    //0x00000de0
        32'h00000000,    //0x00000de4
        32'h00000000,    //0x00000de8
        32'h00000000,    //0x00000dec
        32'h00000000,    //0x00000df0
        32'h00000000,    //0x00000df4
        32'h00000000,    //0x00000df8
        32'h00000000,    //0x00000dfc
        32'h00000000,    //0x00000e00
        32'h00000000,    //0x00000e04
        32'h00000000,    //0x00000e08
        32'h00000000,    //0x00000e0c
        32'h00000000,    //0x00000e10
        32'h00000000,    //0x00000e14
        32'h00000000,    //0x00000e18
        32'h00000000,    //0x00000e1c
        32'h00000000,    //0x00000e20
        32'h00000000,    //0x00000e24
        32'h00000000,    //0x00000e28
        32'h00000000,    //0x00000e2c
        32'h00000000,    //0x00000e30
        32'h00000000,    //0x00000e34
        32'h00000000,    //0x00000e38
        32'h00000000,    //0x00000e3c
        32'h00000000,    //0x00000e40
        32'h00000000,    //0x00000e44
        32'h00000000,    //0x00000e48
        32'h00000000,    //0x00000e4c
        32'h00000000,    //0x00000e50
        32'h00000000,    //0x00000e54
        32'h00000000,    //0x00000e58
        32'h00000000,    //0x00000e5c
        32'h00000000,    //0x00000e60
        32'h00000000,    //0x00000e64
        32'h00000000,    //0x00000e68
        32'h00000000,    //0x00000e6c
        32'h00000000,    //0x00000e70
        32'h00000000,    //0x00000e74
        32'h00000000,    //0x00000e78
        32'h00000000,    //0x00000e7c
        32'h00000000,    //0x00000e80
        32'h00000000,    //0x00000e84
        32'h00000000,    //0x00000e88
        32'h00000000,    //0x00000e8c
        32'h00000000,    //0x00000e90
        32'h00000000,    //0x00000e94
        32'h00000000,    //0x00000e98
        32'h00000000,    //0x00000e9c
        32'h00000000,    //0x00000ea0
        32'h00000000,    //0x00000ea4
        32'h00000000,    //0x00000ea8
        32'h00000000,    //0x00000eac
        32'h00000000,    //0x00000eb0
        32'h00000000,    //0x00000eb4
        32'h00000000,    //0x00000eb8
        32'h00000000,    //0x00000ebc
        32'h00000000,    //0x00000ec0
        32'h00000000,    //0x00000ec4
        32'h00000000,    //0x00000ec8
        32'h00000000,    //0x00000ecc
        32'h00000000,    //0x00000ed0
        32'h00000000,    //0x00000ed4
        32'h00000000,    //0x00000ed8
        32'h00000000,    //0x00000edc
        32'h00000000,    //0x00000ee0
        32'h00000000,    //0x00000ee4
        32'h00000000,    //0x00000ee8
        32'h00000000,    //0x00000eec
        32'h00000000,    //0x00000ef0
        32'h00000000,    //0x00000ef4
        32'h00000000,    //0x00000ef8
        32'h00000000,    //0x00000efc
        32'h00000000,    //0x00000f00
        32'h00000000,    //0x00000f04
        32'h00000000,    //0x00000f08
        32'h00000000,    //0x00000f0c
        32'h00000000,    //0x00000f10
        32'h00000000,    //0x00000f14
        32'h00000000,    //0x00000f18
        32'h00000000,    //0x00000f1c
        32'h00000000,    //0x00000f20
        32'h00000000,    //0x00000f24
        32'h00000000,    //0x00000f28
        32'h00000000,    //0x00000f2c
        32'h00000000,    //0x00000f30
        32'h00000000,    //0x00000f34
        32'h00000000,    //0x00000f38
        32'h00000000,    //0x00000f3c
        32'h00000000,    //0x00000f40
        32'h00000000,    //0x00000f44
        32'h00000000,    //0x00000f48
        32'h00000000,    //0x00000f4c
        32'h00000000,    //0x00000f50
        32'h00000000,    //0x00000f54
        32'h00000000,    //0x00000f58
        32'h00000000,    //0x00000f5c
        32'h00000000,    //0x00000f60
        32'h00000000,    //0x00000f64
        32'h00000000,    //0x00000f68
        32'h00000000,    //0x00000f6c
        32'h00000000,    //0x00000f70
        32'h00000000,    //0x00000f74
        32'h00000000,    //0x00000f78
        32'h00000000,    //0x00000f7c
        32'h00000000,    //0x00000f80
        32'h00000000,    //0x00000f84
        32'h00000000,    //0x00000f88
        32'h00000000,    //0x00000f8c
        32'h00000000,    //0x00000f90
        32'h00000000,    //0x00000f94
        32'h00000000,    //0x00000f98
        32'h00000000,    //0x00000f9c
        32'h00000000,    //0x00000fa0
        32'h00000000,    //0x00000fa4
        32'h00000000,    //0x00000fa8
        32'h00000000,    //0x00000fac
        32'h00000000,    //0x00000fb0
        32'h00000000,    //0x00000fb4
        32'h00000000,    //0x00000fb8
        32'h00000000,    //0x00000fbc
        32'h00000000,    //0x00000fc0
        32'h00000000,    //0x00000fc4
        32'h00000000,    //0x00000fc8
        32'h00000000,    //0x00000fcc
        32'h00000000,    //0x00000fd0
        32'h00000000,    //0x00000fd4
        32'h00000000,    //0x00000fd8
        32'h00000000,    //0x00000fdc
        32'h00000000,    //0x00000fe0
        32'h00000000,    //0x00000fe4
        32'h00000000,    //0x00000fe8
        32'h00000000,    //0x00000fec
        32'h00000000,    //0x00000ff0
        32'h00000000,    //0x00000ff4
        32'h00000000,    //0x00000ff8
        32'h00000000,    //0x00000ffc
        32'h00000000,    //0x00001000
        32'h00000000,    //0x00001004
        32'h00000000,    //0x00001008
        32'h00000000,    //0x0000100c
        32'h00000000,    //0x00001010
        32'h00000000,    //0x00001014
        32'h00000000,    //0x00001018
        32'h00000000,    //0x0000101c
        32'h00000000,    //0x00001020
        32'h00000000,    //0x00001024
        32'h00000000,    //0x00001028
        32'h00000000,    //0x0000102c
        32'h00000000,    //0x00001030
        32'h00000000,    //0x00001034
        32'h00000000,    //0x00001038
        32'h00000000,    //0x0000103c
        32'h00000000,    //0x00001040
        32'h00000000,    //0x00001044
        32'h00000000,    //0x00001048
        32'h00000000,    //0x0000104c
        32'h00000000,    //0x00001050
        32'h00000000,    //0x00001054
        32'h00000000,    //0x00001058
        32'h00000000,    //0x0000105c
        32'h00000000,    //0x00001060
        32'h00000000,    //0x00001064
        32'h00000000,    //0x00001068
        32'h00000000,    //0x0000106c
        32'h00000000,    //0x00001070
        32'h00000000,    //0x00001074
        32'h00000000,    //0x00001078
        32'h00000000,    //0x0000107c
        32'h00000000,    //0x00001080
        32'h00000000,    //0x00001084
        32'h00000000,    //0x00001088
        32'h00000000,    //0x0000108c
        32'h00000000,    //0x00001090
        32'h00000000,    //0x00001094
        32'h00000000,    //0x00001098
        32'h00000000,    //0x0000109c
        32'h00000000,    //0x000010a0
        32'h00000000,    //0x000010a4
        32'h00000000,    //0x000010a8
        32'h00000000,    //0x000010ac
        32'h00000000,    //0x000010b0
        32'h00000000,    //0x000010b4
        32'h00000000,    //0x000010b8
        32'h00000000,    //0x000010bc
        32'h00000000,    //0x000010c0
        32'h00000000,    //0x000010c4
        32'h00000000,    //0x000010c8
        32'h00000000,    //0x000010cc
        32'h00000000,    //0x000010d0
        32'h00000000,    //0x000010d4
        32'h00000000,    //0x000010d8
        32'h00000000,    //0x000010dc
        32'h00000000,    //0x000010e0
        32'h00000000,    //0x000010e4
        32'h00000000,    //0x000010e8
        32'h00000000,    //0x000010ec
        32'h00000000,    //0x000010f0
        32'h00000000,    //0x000010f4
        32'h00000000,    //0x000010f8
        32'h00000000,    //0x000010fc
        32'h00000000,    //0x00001100
        32'h00000000,    //0x00001104
        32'h00000000,    //0x00001108
        32'h00000000,    //0x0000110c
        32'h00000000,    //0x00001110
        32'h00000000,    //0x00001114
        32'h00000000,    //0x00001118
        32'h00000000,    //0x0000111c
        32'h00000000,    //0x00001120
        32'h00000000,    //0x00001124
        32'h00000000,    //0x00001128
        32'h00000000,    //0x0000112c
        32'h00000000,    //0x00001130
        32'h00000000,    //0x00001134
        32'h00000000,    //0x00001138
        32'h00000000,    //0x0000113c
        32'h00000000,    //0x00001140
        32'h00000000,    //0x00001144
        32'h00000000,    //0x00001148
        32'h00000000,    //0x0000114c
        32'h00000000,    //0x00001150
        32'h00000000,    //0x00001154
        32'h00000000,    //0x00001158
        32'h00000000,    //0x0000115c
        32'h00000000,    //0x00001160
        32'h00000000,    //0x00001164
        32'h00000000,    //0x00001168
        32'h00000000,    //0x0000116c
        32'h00000000,    //0x00001170
        32'h00000000,    //0x00001174
        32'h00000000,    //0x00001178
        32'h00000000,    //0x0000117c
        32'h00000000,    //0x00001180
        32'h00000000,    //0x00001184
        32'h00000000,    //0x00001188
        32'h00000000,    //0x0000118c
        32'h00000000,    //0x00001190
        32'h00000000,    //0x00001194
        32'h00000000,    //0x00001198
        32'h00000000,    //0x0000119c
        32'h00000000,    //0x000011a0
        32'h00000000,    //0x000011a4
        32'h00000000,    //0x000011a8
        32'h00000000,    //0x000011ac
        32'h00000000,    //0x000011b0
        32'h00000000,    //0x000011b4
        32'h00000000,    //0x000011b8
        32'h00000000,    //0x000011bc
        32'h00000000,    //0x000011c0
        32'h00000000,    //0x000011c4
        32'h00000000,    //0x000011c8
        32'h00000000,    //0x000011cc
        32'h00000000,    //0x000011d0
        32'h00000000,    //0x000011d4
        32'h00000000,    //0x000011d8
        32'h00000000,    //0x000011dc
        32'h00000000,    //0x000011e0
        32'h00000000,    //0x000011e4
        32'h00000000,    //0x000011e8
        32'h00000000,    //0x000011ec
        32'h00000000,    //0x000011f0
        32'h00000000,    //0x000011f4
        32'h00000000,    //0x000011f8
        32'h00000000,    //0x000011fc
        32'h00000000,    //0x00001200
        32'h00000000,    //0x00001204
        32'h00000000,    //0x00001208
        32'h00000000,    //0x0000120c
        32'h00000000,    //0x00001210
        32'h00000000,    //0x00001214
        32'h00000000,    //0x00001218
        32'h00000000,    //0x0000121c
        32'h00000000,    //0x00001220
        32'h00000000,    //0x00001224
        32'h00000000,    //0x00001228
        32'h00000000,    //0x0000122c
        32'h00000000,    //0x00001230
        32'h00000000,    //0x00001234
        32'h00000000,    //0x00001238
        32'h00000000,    //0x0000123c
        32'h00000000,    //0x00001240
        32'h00000000,    //0x00001244
        32'h00000000,    //0x00001248
        32'h00000000,    //0x0000124c
        32'h00000000,    //0x00001250
        32'h00000000,    //0x00001254
        32'h00000000,    //0x00001258
        32'h00000000,    //0x0000125c
        32'h00000000,    //0x00001260
        32'h00000000,    //0x00001264
        32'h00000000,    //0x00001268
        32'h0ff000ff,    //0x0000126c
        32'h00000000,    //0x00001270
        32'h00000000,    //0x00001274
        32'h00000000,    //0x00001278
        32'h00000000,    //0x0000127c
        32'h00000000,    //0x00001280
        32'h00000000,    //0x00001284
        32'h00000000,    //0x00001288
        32'h00000000,    //0x0000128c
        32'h00000000,    //0x00001290
        32'h00000000,    //0x00001294
        32'h00000000,    //0x00001298
        32'h00000000,    //0x0000129c
        32'h00000000,    //0x000012a0
        32'h00000000,    //0x000012a4
        32'h00000000,    //0x000012a8
        32'h00000000,    //0x000012ac
        32'h00000000,    //0x000012b0
        32'h00000000,    //0x000012b4
        32'h00000000,    //0x000012b8
        32'h00000000,    //0x000012bc
        32'h00000000,    //0x000012c0
        32'h00000000,    //0x000012c4
        32'h00000000,    //0x000012c8
        32'h00000000,    //0x000012cc
        32'h00000000     //0x000012d0
    };
    
    logic [11:0] instr_index;
    logic [31:0] data;
    
    assign instr_index = i_addr[13:2];
    assign data = (instr_index>=INSTR_CNT) ? 0 : instr_rom_cell[instr_index];
    
    always @ (posedge clk or negedge rst_n)
        if(~rst_n)
            o_data <= 0;
        else
            o_data <= data;

endmodule
